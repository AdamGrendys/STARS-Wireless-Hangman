/* UART Transmitter File
Descriuption: x
*/

module uart_tx (
    input logic clk, nRst
);


endmodule