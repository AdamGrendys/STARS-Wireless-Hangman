/* TLCD Controller (Provided)
Descriuption: x
*/

module lcd_controller (
    input logic clk, nRst
);


endmodule