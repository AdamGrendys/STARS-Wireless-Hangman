/* Keypad Controller for Host File
Descriuption: x
*/

module keypad_controller_host (
    input logic clk, nRst
);


endmodule