/* Top File
Descriuption: x
*/

module display_fsm (



);


endmodule