/* Top File
Descriuption: x
*/

module main (



);


endmodule