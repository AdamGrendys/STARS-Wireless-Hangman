/* Top File
Descriuption: x
*/

module game_logic (



);


endmodule