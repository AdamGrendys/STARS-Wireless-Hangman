/* Host display for game logic
Description: 
*/
