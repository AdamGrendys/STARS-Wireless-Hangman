/* Top File
Descriuption: x
*/

module KeypadControllerPlayer (



);


endmodule