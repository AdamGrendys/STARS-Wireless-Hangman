/* Top File
Descriuption: x
*/

module top (



);


endmodule