/* Top File
Descriuption: x
*/

module keypad_controller_host (



);


endmodule