/* Display FSM File
Descriuption: x
*/

module display_fsm (
    input logic clk, nRst
);


endmodule