/* Top File
Descriuption: x
*/

module buffer (



);


endmodule