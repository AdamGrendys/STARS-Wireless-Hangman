/* Keypad Controller for Player File
Descriuption: x
*/

module keypad_controller_player (
    input logic clk, nRst
);


endmodule