/* Top File
Descriuption: x
*/

module keypad_controller_player (



);


endmodule