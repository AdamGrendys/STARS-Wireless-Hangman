/* Top File
Descriuption: x
*/

module msg_reg (



);


endmodule