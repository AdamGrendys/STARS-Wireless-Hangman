/* Top File
Descriuption: x
*/

module lcd_controller (



);


endmodule