/* Game Logic File
Descriuption: x
*/

module game_logic (
    input logic clk, nRst
);


endmodule