/* Main File
Descriuption: x
*/

module main (



);


endmodule