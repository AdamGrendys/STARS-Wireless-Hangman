/* Top File
Descriuption: x
*/

module uart_rx (



);


endmodule