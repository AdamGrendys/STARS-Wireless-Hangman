/* Top File
Descriuption: x
*/

module KeypadControllerHost (



);


endmodule