/* Message Register File
Descriuption: x
*/

module msg_reg (
    input logic clk, nRst
);


endmodule