/* UART Reciever File
Descriuption: x
*/

module uart_rx (
    input logic clk, nRst
);


endmodule