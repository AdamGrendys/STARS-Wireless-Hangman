/* Top File
Descriuption: x
*/

module uart_tx (



);


endmodule